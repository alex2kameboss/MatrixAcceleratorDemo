`ifndef CVA6_PARAMETERS_SVH
`define CVA6_PARAMETERS_SVH

// AXI parameters
`define CVA6_AXI_ADDR_WIDTH 64
`define CVA6_AXI_DATA_WIDTH 32
`define CVA6_AXI_ID_WIDTH 4
`define CVA6_AXI_DATA_USER_WIDTH 1

`endif // CVA6_PARAMETERS_SVH