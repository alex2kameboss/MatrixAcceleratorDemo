module matrix_accelerator_subsystem (
    input   clk     ,
    input   rst_n   
);
    
endmodule