`include "soc_parameters.svh"
`include "axi/typedef.svh"

module matrix_accelerator_soc (
    input           clk     ,
    input           rst_n   ,
    output          tx      ,
    input           rx      
);

typedef enum int unsigned {
    RAM             ,
    UART            ,
    AXI_NO_SLAVES   
} axi_slaves_e;

// Local Parameters -----------------------------------------------------------
localparam AXI_NO_MASTERS = 2;

localparam AXI_DATA_WIDTH   = `SOC_AXI_DATA_WIDTH;
localparam AXI_STROBE_WIDTH = AXI_DATA_WIDTH / 8;
localparam AXI_ADDR_WIDTH   = `SOC_AXI_ADDR_WIDTH;
localparam AXI_USER_WIDTH   = `SOC_AXI_USER_WIDTH;
localparam AXI_ID_WIDTH     = `SOC_AXI_ID_WIDTH;
localparam AXI_ID_WIDTH_SLAVE = AXI_ID_WIDTH + $clog2(AXI_NO_MASTERS);

localparam RAM_LENGTH = `SOC_RAM_LENGTH;
localparam RAM_WORDS = RAM_LENGTH / AXI_STROBE_WIDTH;

localparam UART_LENGTH = 2 ** 5;

localparam axi_pkg::xbar_cfg_t xbar_cfg = '{
    NoSlvPorts:         AXI_NO_MASTERS,
    NoMstPorts:         AXI_NO_SLAVES,
    MaxMstTrans:        4,
    MaxSlvTrans:        4,
    FallThrough:        1'b0,
    LatencyMode:        axi_pkg::CUT_MST_PORTS,
    PipelineStages:     0,
    AxiIdWidthSlvPorts: AXI_ID_WIDTH,
    AxiIdUsedSlvPorts:  AXI_ID_WIDTH_SLAVE,
    UniqueIds:          1'b0,
    AxiAddrWidth:       AXI_ADDR_WIDTH,
    AxiDataWidth:       AXI_DATA_WIDTH,
    NoAddrRules:        AXI_NO_SLAVES
};


// Data Types Definition ------------------------------------------------------
typedef logic [AXI_DATA_WIDTH-1:0] axi_data_t;
typedef logic [AXI_STROBE_WIDTH-1:0] axi_strobe_t;
typedef logic [AXI_ADDR_WIDTH-1:0] axi_addr_t;
typedef logic [AXI_ID_WIDTH-1:0] axi_master_id_t;
typedef logic [AXI_ID_WIDTH_SLAVE-1:0] axi_slave_id_t;
typedef logic [AXI_USER_WIDTH-1:0] axi_user_t;

`AXI_TYPEDEF_ALL(master_axi, axi_addr_t, axi_master_id_t, axi_data_t, axi_strobe_t, axi_user_t)
`AXI_TYPEDEF_ALL(slave_axi, axi_addr_t, axi_slave_id_t, axi_data_t, axi_strobe_t, axi_user_t)

typedef enum logic [31:0] {
    RAM_BASE  = `SOC_RAM_BASE   ,
    UART_BASE = `SOC_UART_BASE   
} soc_bus_start_e;


// Wires ----------------------------------------------------------------------
logic                               ram_req;
logic                               ram_we;
logic [AXI_ADDR_WIDTH - 1 : 0]      ram_addr;
logic [AXI_DATA_WIDTH / 8 - 1 : 0]  ram_be;
logic [AXI_DATA_WIDTH - 1 : 0]      ram_wdata;
logic [AXI_DATA_WIDTH - 1 : 0]      ram_rdata;
logic                               ram_rvalid;

AXI_BUS #(
    .AXI_ADDR_WIDTH ( AXI_ADDR_WIDTH    ),
    .AXI_DATA_WIDTH ( AXI_DATA_WIDTH    ),
    .AXI_ID_WIDTH   ( AXI_ID_WIDTH      ),
    .AXI_USER_WIDTH ( AXI_USER_WIDTH    )
) master [AXI_NO_MASTERS-1:0] ();
AXI_BUS #(
    .AXI_ADDR_WIDTH ( AXI_ADDR_WIDTH        ),
    .AXI_DATA_WIDTH ( AXI_DATA_WIDTH        ),
    .AXI_ID_WIDTH   ( AXI_ID_WIDTH_SLAVE    ),
    .AXI_USER_WIDTH ( AXI_USER_WIDTH        )
) slave [AXI_NO_SLAVES-1:0] ();
axi_pkg::xbar_rule_32_t [AXI_NO_SLAVES - 1 : 0] routing_rules;

AXI_LITE #(
  .AXI_ADDR_WIDTH   ( AXI_ADDR_WIDTH ),
  .AXI_DATA_WIDTH   ( AXI_DATA_WIDTH )
) axi_uart ();


// Combinatorial Logic --------------------------------------------------------
assign routing_rules = '{
    '{idx: RAM , start_addr: RAM_BASE , end_addr: RAM_BASE + RAM_LENGTH  },
    '{idx: UART, start_addr: UART_BASE, end_addr: UART_BASE + UART_LENGTH}
};


// Modules Instantiation ------------------------------------------------------
matrix_accelerator_subsystem  i_core (
    .clk         ( clk      ),
    .rst_n       ( rst_n    ),
    .boot_addr   ( RAM_BASE ),
    .core_axi    ( master[0]),
    .acc_axi     ( master[1])
);

// axi interconnect
axi_xbar_intf #(
    .AXI_USER_WIDTH ( AXI_USER_WIDTH            ),
    .Cfg            ( xbar_cfg                  ),
    .rule_t         ( axi_pkg::xbar_rule_32_t   )
) i_xbar_dut (
    .clk_i                  ( clk           ),
    .rst_ni                 ( rst_n         ),
    .test_i                 ( 1'b0          ),
    .slv_ports              ( master        ),
    .mst_ports              ( slave         ),
    .addr_map_i             ( routing_rules ),
    .en_default_mst_port_i  ( '0            ),
    .default_mst_port_i     ( '0            )
);

// memory
axi_to_mem_intf #(
    .ADDR_WIDTH ( AXI_ADDR_WIDTH    ),
    .DATA_WIDTH ( AXI_DATA_WIDTH    ),
    .ID_WIDTH   ( AXI_ID_WIDTH_SLAVE),
    .USER_WIDTH ( AXI_USER_WIDTH    ),
    .NUM_BANKS  ( 1                 )
) i_axi_to_mem (
    .clk_i          ( clk           ),
    .rst_ni         ( rst_n         ),
    .slv            ( slave[RAM]    ),
    .mem_req_o      ( ram_req       ),
    .mem_gnt_i      ( ram_req       ),
    .mem_addr_o     ( ram_addr      ),
    .mem_wdata_o    ( ram_wdata     ),
    .mem_strb_o     ( ram_be        ),
    .mem_we_o       ( ram_we        ),
    .mem_rvalid_i   ( ram_rvalid    ),
    .mem_rdata_i    ( ram_rdata     ),
    .busy_o         ( /* Unused */  ),
    .mem_atop_o     ( /* Unused */  )
);

tc_sram #(
    .NumWords   ( RAM_WORDS         ),
    .NumPorts   ( 1                 ),
    .DataWidth  ( AXI_DATA_WIDTH    ),
    .SimInit    ( "random"          )
) i_dram (
    .clk_i  (clk_i                                                                          ),
    .rst_ni (rst_ni                                                                         ),
    .req_i  (ram_req                                                                        ),
    .we_i   (ram_we                                                                         ),
    .addr_i (ram_addr[$clog2(RAM_WORDS)-1+$clog2(AXI_DATA_WIDTH/8):$clog2(AXI_DATA_WIDTH/8)]),
    .wdata_i(ram_wdata                                                                      ),
    .be_i   (ram_be                                                                         ),
    .rdata_o(ram_rdata                                                                      )
);

// uart

axi_to_axi_lite_intf #(
    .AXI_ADDR_WIDTH     ( AXI_ADDR_WIDTH    ),
    .AXI_DATA_WIDTH     ( AXI_DATA_WIDTH    ),
    .AXI_ID_WIDTH       ( AXI_ID_WIDTH_SLAVE),
    .AXI_USER_WIDTH     ( AXI_USER_WIDTH    ),
    .AXI_MAX_WRITE_TXNS ( 1                 ),
    .AXI_MAX_READ_TXNS  ( 1                 ),
    .FALL_THROUGH       ( 1'b0              )
) i_uart_axi_to_lite (
    .clk_i      ( clk ),
    .rst_ni     ( rst_n ),
    .testmode_i ( '0 ),
    .slv        ( slave[UART] ),
    .mst        ( axi_uart )
);

uart_mock i_uart (
    .clk    ( clk       ),
    .rst_n  ( rst_n     ),
    .axi    ( axi_uart  ),
    .tx     ( tx        ),
    .rx     ( rx        )
);

endmodule